module acpi