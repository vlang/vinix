module sys

pub const (
	KERNEL_VERSION = "0.1.0"
)