module memory

const page_size = 0x1000
