module main

fn main() {
	println('fetch placeholder')
}
