module sys

pub struct Mutex {

}

pub fn (mutex &Mutex) lock() {
	//TODO Implement mutex locking
}
