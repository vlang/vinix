module sys

