module time

pub struct TimeSpec {
pub mut:
	tv_sec  i64
	tv_nsec i64
}
