module sys

const (
	kernel_version = "0.1.0"
)