module public

pub const af_inet = 1

pub const af_inet6 = 2

pub const af_unix = 3

pub const af_local = 3

pub const af_unspec = 4

pub const af_netlink = 5

pub const sock_nonblock = 0x10000

pub const sock_cloexec = 0x20000
