module memory

__global ( page_size = u64(0x1000))

__global ( higher_half = u64(0xffff800000000000))
