[manualfree] module errno

pub fn get() u64 {
	return 0
}
