module main

import os

fn main() {
	println('Vinix Init started')

	for {
		os.system('cd ~ && bash --login')
	}
}
