module sys

pub struct Mutex {

}

pub fn (mutex &Mutex) lock() {
	
}