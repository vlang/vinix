module sys

const (
	KERNEL_VERSION = "0.1.0"
)