module acpi

fn lol() {
	
}