module main

fn main() {
	println('mount placeholder')
}
