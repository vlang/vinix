module sys

pub fn (kernel &VKernel) get_cmdline_option(name string) string {
	return ''
}